BZh91AY&SY�W;P -߀Pxg����߰����P>:m��8Z���$�Ѡ�F�'�ďɡ���P��@�=&��hh �   �#PI�@ё��    2d�b`ɂd ф``"	��i�G�f����=C#C���i ���IU�D Eш4%(O��_�h�Va �7�g�	�tc<�*��* 1�b�G�� ��g�OA��rb?~4�O��K���A|xS[x#g�wg�+���d`�K��ph�5:���rGVIRs��n��G��<L�0�p�<$
�T���u�2w�L�]a����ׄU��2���v;3&M7gkW&[�U�p71Ƚ&���jN�9�pP�$@�A�D�"�5�y�B,?d.�����48{D�U��;����<D�(�S"��.鴄ecF
��V�BF�Z��3`cH�U��agV.�J��s�5��calZ44�z(f�W=�^0��|��-����m��A���?���$�|
OH���@��"
�G�a?[@6)nȁ�IK�(U�j"b��NfjZ�jռ����f���ǳ��K<��mn�k�ڗe����{}�_%&2xg�u�DfZ���𞅂�����~2�W.�	jZ!|�N�7-ҷa���f~�3$���-%F�ϬɅ(�zg��4q#Ǜ�c)�`^w�t����󬇷q�-�62�R@�)�µ�IsP3�7�K���2�!T2��4-�]��Rj'��
A�0~�~F4�Af�	��s
�������3�
0?`������`_Yi\c<9����T͖�eRu��(� �Ί� 
����.�K��j�"��f2H�����X����&��&Ӗ����X�3'ʠjf��p>��*030�a�E�_�ƞ63O���M�^���� +u�q`rZ�lm�2� 4F����1r�V�r
"I#IJ�]��:K�Q-�ZG���3��T���w/)�4U(VѠ+
�yb�Ju��x�n�l�K�Z�I��#��������4ϒ�o�Y7z��̵����]�1^�� N�n�R�7*q9r��r�I0�!)��S ��u��iJ�aA��|�����9�V�R丬�g3E���a�r�?5H��IK�Y%1G���6�F�Q
��r{�&FH�A�f��*)�]П8�&N�dD�;ށ�S���2�!��[�.)�m�C*�
��\;]�EˑPI�����A�� �OD�Q/�]��BCy\�@