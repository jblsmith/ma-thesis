BZh91AY&SY`�̏ �_�Py����߰����`�y�N!�aݔ 8J�i4�zQ��H   �ј�P��2@     ��!�	�4ѣ4ɑ� �DB
i�MCM�i�OSF�26H  i��ɂ0�#M1L� $�@���y���A=&�dyC�@�ԺI&�|���.�$Y�O��ր�A�Π�g���h/_�K�������>�p(��@�bY��d�\�
����A��94�Y}�2�͙�E\���eb��z�k-�1}bIg�ApUC��C��jk�V
a���C#�]�2����;�hc$� �j֣eZ�p�H 7w�ݱƂ9Ǎ�2�\�|���-�VZV���.��ɷv_�6�;�@�Q�,���k�oSm�Ԛz�z���b��QS\``��CN���x�N[n4�SyS{r-כ-љ�}����5-�H0����|A�9+d�)�(�O �"����td3�M�i��5�gycw�b����Asmk"���(TqkP<�d{�d����)���
��֥WZ(�0A+��nZMJD3f��9#�n�qu{w,f��v�qX��JRJ��d��VZh�UF(�ҫ=��#UC�8X���ܖR��P�����������L�ccT���2��0����C.[~s�s�I�61���m�ؚBPAC��HI�l�*),T���$���e$�s0W�E��%i��!��9���pp��JG+%+C�i�R�̔����\�N�&MtD��������q�òh�$1�M���@�̓gu�j�#�}e�H�Q�@�l�4��K&�'��o�d��h�#(��0��ҙ7NڎL����zOG���rS������h�T$�YJ���{$}�l�V������̥�NՒ���ܻ�5;�?/��}𓄟8����Խ�L��ϫ7���a�ݶ-(Yc�����a��#lU1���8S�V���#�7��?��i�Y�D)�/�t�G��5G���/��U�dtੑ��ޤb��M8ʔ�2b����f+#r2|B�!.����PT�Qc��y�.d�Ǒ��4s�1[����s����9'�����t_�i��S�pU��Ҷoǧ�t$ѵJ�Eof���ϰ�\��˝W�S�Y��.���+HI�y�cr��k��uɢ��e�6.�ɋf1�oa�.R�v%ȅ)h�o�����t�vU��S��c�6�V*\IFE	D�"Z,aT$�(�wO���I]�lNp���b>g\�7���{~L��j?���o.��:us�|�qآS�SœeH�͂�BJtaz�^�T���X��=.������k��[7c��Q�x14�h�R��e�u��0q�3�av�꽺~,�k�f�h���-^�zi�_���f4�N����x����q���\���1���*�Mʜ&Q�v�k�6��v�ۜ���$ǈ֝_:�Y��7/����M������u�c��}T�/��ɣ��Y'j����y�,#�rE8P�`�̏