BZh91AY&SY7k'V ߀py����߰����P���`�k�2�i�$�@L?MOL�BdA�� �� 4�OBQ�=M<��2  DDLL���6�!��i�&OP ��i��ɂ0�#M1L� $H@�D���SП�~�SCjM24  !Tk�d!�H�	��Н�=��j?�
��l[��K�=��m* _� 1�yZ��Ʈ~L�7]��>d����}��F��������(A�ǯtuM��EE������b�n�8�#z���~�s�Y{$fs�d]�ƾ�4(4�������G�������9�pqن]|�����bCi�^.��yd�:c#8�3S8;m��z�JA�x�#��e�!�хi�-M� �)`���޺��i�|�W|���rZ(�H���"q�9�^/J!kTBִE�(��EMd���$L��QT�5����B�:λ�K��]�@.���x7j�0�$�F���`�DS���R�y���߈������,����c5�B��	jR��EX5
b�Л�XԵ^��4����\���I�ۏ���O�3�/n��>�d=G��\�͟��M^+�VT�ޢ��w���H��}���Oؗ_n&�#���?U�ֻ_����hF�c-����|�#�H�ɞK{���q3�H%�>1#�2{*!`i,7b^	�
wvN���	�&��o&
^�Ճ+JJ�����6bkCV:�������� i*`@%��jwH��&b崍E�bl�!ťe�����1J������=���v��+	g��GTѽK�'2Ng����KԎ���[�BEwR�8�Ġ��)w9!��m�8jk��F�H�>�fj�g��D{)Mf�j��ߔ 
	T�p�4�O�MP/�4żJ+EN�Q<��"���щ`WD��Y#��@͐�A��T��Kd��J�l�j�YP*��|zD=�U�8ȋ]�h{�� ���U@th[�֜-�0�ٺ6��3�j2�*��$X������%�˔��6j����Ҕ�]��
de"�a����[����:�A�:�1}��b�e����\�a���1��� ���c�'�xX��d�"�b�E]4�8[�4���b���G�(#h�Yt%�lZ�������V]��fX(I���;�x2���O�]��B@ݬ�X