BZh91AY&SY�� ~_�px���������`?ݹ`���(�]�$�b�d	�5���&���Cdz�4�@��h�h      q�&�a22bh�A�L 4���Q��M4�M��L 4� q�&�a22bh�A�L $DF��#SSM�<Sb	�h���`� K#�BX1"@B H��JD�п��Z����X6��}l�TaI�~Z�!�o�Y������]����k�ӭ���Ϯ�����à��̂��k�ܚ<$�t�g�0�d���)s���L��u�B�˱�F�ݷP��b-dX�4]l'5��3	�D��
�l!��Q=:Fk,ժ*�r�%R�$�p�=!���,����Y�篧��r!6�ӥx7��-Q�8w�8I����[�����)B���vv��	�t)l�X��,ս���$CA�2�a�A��%�	Pƶ�F�R�VR�bFMN�=�#SeEb↹�j�ɋ,�2��A��˺�* ;]��6:0a�=-�qLe6!Sa�o��f"�儊��2(K�[J	,�&��Վ�b��-)�ś�ah��E!���:`�f�MV���+R��$FـN;�87ӮVES;0q�m�l���eN�l�X���k�m�� ���P���䷫�%�Dr��U��]7��-��{�C�)�&"$��B�! ��*�!�a�Q��eh�OC��tГ&jZ�1���HWaw��������c�G3�z�:���X�}���Wx1��E�����X�aWu�j�F���������͟���7�%���0��y���ga��F�!{�|8�>/�p��X�hl��1�u�!v��ya��B"�	����w�c{H����V􋒲�mɿ���ڛ"��A�Q
���>h�gZ���Y߳20O\��K;�֍��Z��!�OJpo��)MU��`�!�ƓM:�D����(08�������,)��]a=�
�+)�{��)�,��h(%U6�:���B�Y���[�K��_�g�*HP��E��Ňea`��
�5���0��d�=�n*.5@(.�H�1kk��Mj�M.�sh!f��0�h������&�(K&8��+\-5��0.O���k���*1nv��@����$4��Z*����Ju&�  ,�T䦒P|j�bLdz' ΘGD\X5�T'��G��pQ,�x��B�Po�oe)͍�����$����+�
�b~_y����I��=�d�.�o��3��d��q1�,e����;���\�f`��.�6����(�ef��V�GT�:"���N����S�^pܼ�T`kt����\�����9q%�Kb9c�� �l��=���6B����;��ײ�{H��2�%�Q�Z��v����2~~���c�f�v�XB�dkP��������E�F�ad����)����h