BZh91AY&SYl�a� �_�Py����߰����Px+#i�ۉ�\�IM��=L�i��i�=2�h�hM4d �M Ч�S�?H�# �     ��@JiL���4�#�@2z@q�&LF& L�&@F �$D=M��OPmC� h4  ),�(H�J�"�I�_�ʃ?��X���2Z�~��:��W -cta�Դ�{��9������G3���p���&T�>����H8�q���gèq�E��C�k��|<`�8.������I%Jrȁ^����C�PqQ�m�v�HfL�L�l��D��͎�D�[j��߭�2I��8z&�o�r�҇/�'���E����� ��n���;�Pl���W���DΌ�s`�3W�UWKMp+
�pH_�nmѼ�[cco��l( �%�U>	G��5"�c���몙�m�AXd(-�m��β�A��u����	vaa7��R՛���	E�ڦ=�����E�WX�:��GK}b������Mz<<�ϋ?I�	~�;����B
�f��HT(V��5w<�J�-B�Y�%ܵA��{�"��̑�9�'/Qs�m��6Dx'�؊-r��x���!�	B�i�2��%,L+c $�1nɎ�N0�Yw×&�2 �$�d�F�3-�L��<�R@+6�}��F0,�@&Lj&���3����X�yʧ���c&��Y�Y�1��a��f��NH�Aˌğ�>B�m�A��r?48�F�/',-��P��y1�brp�d}��&d��fa��3b��*x޷��^L�p��4R7�-6EC�Y=�lD.�<���+�$Ti���IH��	�u�x�â[�W5Ă@�x_�PZ,��nsR���A5�j�!b*����!���7w�5��!K��\���/��A����
���9���g�9KK&��4Xd���ҭY1u�(WRC��̚Rx��:��
z�+P'�6<6�T�N���*��Y�05�AI���ApZ(��a��z�a����P;�-!i�(1`�[��{�Y1�d9�zס�Ԭ6�pP�����܌�����"̮RK�l��A�� �N��]��BA����