BZh91AY&SY�.M _�Py����߰����`�      T�OI=A���4� �@�bC��2b10d�2 h�00dɓ��&	�F�!��&L��L �0L�0�2d�b`ɂd ф``"	� #M=4�&������H�5�@Th� �E���	H/�/����0��A ��J!K_c���D}K�bY�!\i�/Ь@I+��V�u#0D}��@�T�I���BRCvs0?���4�̳��x��u�J$��ΧP�b�>9Je}gXe"��,YM��]r���I^E��3i�pI��)���HT.I�3�d#<����&�w��S{�PU�P�+j� �����^O�]�'��<(��gi�z��m0�$�CO��|C:�<�H�4���3���IP�$�gI+V:�cϚ��AB�DQ����Vv�3H!P��$�C�Qj�v�y�q*�E9J��rL�F�I&&lAWK�"�۶���1�20�It�Q��J��B��u-%���f�b���*L��rC2r�xR5B�3��\x�r-%����3.`��rT�P��c6�c+�2�w1A�t��!�R�6ɝ2��V��5dj��h�S3:K�<T���Vz(f�_H��:�<�����o��m�1$�����$�H��TRX����T}��a}�h�(^	(_�?�Y����`P��%$T`0��LT̠I���	j����`��N�������W�?S7撗�<Q���C�����}�����ڴ���c���a�Ӕ������V �>)��t
�X��.�Ƈi�c��h��Q$��e�_����ǂ]f1�I�F1��	+Z��~	�I�qo����d@�T�T�����B?~��zp$�	v��clcc����C�fILʦ�נ+��H���p�%�{�,�q���/x+�~��;��8�eko�%�F����PcEX`����0j�%h�����0*4��	'��W�t����G����)�����\UFE�kG���K�쐹�s[�@0IPtvC��D�9���sw {K�7zL��Ƹ�K�q�`8NB��p����3pBzl�Ҧ��	,�6�=�C'����xy��r����J6��!@����g�>�aD�2C� ��9I$��\�*l�����(Hd#۵Y#�(��*Ħ`  �̀�*��#@�U�*\���X�h�{�@_���}��8�%�T�i��s�P_��c�X��5�������d���&P;YsSH�A�	&q�t:�� Ν�s�`��u�0�̍�!��0�����
�5�A.�yT��*�TH�k^G n'z�(d5��}_%Ac��6����f^��r��Kv�����i�N��8����5�5�Y���0-F�#�JW�T+�h�>$���`q����cZ���o.]�.]��5KP�x�c�@���p��ۥ����)�w�rh