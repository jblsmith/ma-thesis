BZh91AY&SY�>2� D߀py����߰����P�qGエ@�#L�)�OM&����� ɓ@=&�2J �      a�������@� �� d4��d�L����L� $&�h�di���4�  4�L�I+�hƄI	""�{�$'�H��3C��V��gZBra�.���h��6 �#b-*��P��͇K�|���ۘ�s
"]t<z\?�̙�ժ����[�6Yڊ�N��e�Q�|:R}���d
��^<1��H�3��E7�$�
W	�t�h����G&�Ggo�sˀD��EOw57��^���� w <���B��H� F����X� +4ݹ� 	B���q ڄ]l	�y���P*!���lr���Ϣ�k�5�]`�W=����hrYEe3H0�H�B2������*��j��5� X�T*����	p�j�hU�5��Ԡ�NH�Q'_���9�}���,� @P@ 	a��g�D�h�wە��h�H��2yQ2:�^%!CA�X)D� �$Y�K�"�Q�iÕ��'.�1Z�ϖQ�J4���h�O:��z��]����_׮ҵ�����j��xS�ꢻ�;f~�Ǎqѷ��@Tg�+?�}�|[����1����'/�v�s��ƜD��h�4uӻ�3P�f�[9��9��Q��ʢP��|t�-Ć�BѴ\���G. WMF+,���8;6²�*21*�,��8���
	o����)����,���ɰ>�	��MZR�o%`�tav�ǕT��ʪ+G�,mG���i�08!M2r��zҟa�C>�0�8�P��(��f}F3D��R�P̯B���d��Z�fa���}�3(����+�Ӻă2B��"����|jap�i��CrH���	�y*I
�m�~&tL��q	�����DE�L��$M��D�j�!D%	�"���Ǻ!�6T�a���R�>3Kl��珘�:6Q���a^��h9�3*���H���	��mL=��dw�'.N��M����6��T#�"���Pa��õ]�4�ɟ:{>ç�L�&b�#O��Q�`���¸4g��iD j�;�cA!J��s7����*�������.�T`;4�6BHr'��\*���$�]^�9��V�ܦ�ܟ����4>�)9w9fL����d��]��BCD��D