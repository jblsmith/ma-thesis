BZh91AY&SY^X| 
߀Px����߰����P~p��6�l�"���F��	�mS���6�ѩ��=@�l�i��H       " ��Ч�<��z�2<�� 4 �0&&�	�&L�&	���R�z'� �   �5�}��AB@����;܆�'䖨Fl8�H'#ޑ ��l�1�#sR�Y���Y������u�K��H�"�u��sGK+M�-<��x�y�ʝ�4��f2|3N���tfj�h���m�a���Qj�T����ג	x49��4�ƑT��2�(��G�0�9�N���xe�Y
Hm4�w��W:�c��dZ/s3gT6�<xo�3��G�r3[b�0��<m��S��3Xn7AǑ�3���|c�J[+)�2xD��^!����#:��u
�e�5�(]i��1��A�����z��[)�X����^)Yp��P�
��������)ddXF�N':�fb\e�.$15�Mq���&�Y֖�
vd��B�S�7$.��e[��8�.Erܡj������;M����m�A��<%��	�R'lRl�>[)�,0��^Y @����;�@�*�IK��$`��
b�J�����̽��^��k�|a�\�e]~Ʋ��] ���l�������^XS-ޭ�%��ٟ��S]��L@��:��~q&I@�_ˤN�d��2@/��GƊ�m/�<��ֈ�S��B���2�f4�M���Ċ�ɢ]+�5��Fl��.]�$v�P�롶�nc��iT)�1����ڂ�����m`��F6�d�~񫚇3OJ�t�2D��i���Z��T"z�4�e�8ᕴ�V\) z*��6ig5I,qJC�z�=�*с%I9�����#�ql��I"���D�-�yo�Z�^Jr~�(ra���VҳQ��#���2����:�F��*-m����}pQtc���m�Ho*�FѸ6IuJ�#jp�+�����b�J+EMD@�RRavBӘ�z%�%�P�!8L�ePgU[��T؝�S���- 2h�տxH����r��D\4�4��8zwQШ<&��W�-_vѰ��w���V�Jv4�3����P"��@p�$�*h�r%#N�jT��
��DX��ߠ�!)�抙�{�Χ�^j�[�6�����.+.-��27OL���9B��%`�O]�轐V2�}�UPi�*���QG���ko���˼b߿ه�n�ì�d`n��Kk5=|����A-4ퟞ�e���"�(H/�> 