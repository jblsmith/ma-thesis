BZh91AY&SYP�� Y߀Py����߰����P�n�wc��閐ILh4�4d�OS����i�P��4LF��C�hz�� M&�H��B�Q�Q����A��2d�b`ɂd ф``I2M��L&��&�  EH3�@�"T�2,T$�uׯ���K\����I��R� ��P��@	 �B�P	)G^�����8��ơ�����E�"x�g���iO��$S�k�Ǟ<1��$t��	P-گ�+�-����h�ɾXQ��2��k�8����@/s��ϝ�P�d�V~�e��8���I�2iq[-[�������pckOe��
�v�f]�m����p�u�gvJ�t�(�����as�`�L"V�$E�_a��B�]�k�H��Co)!�-�elQ�hM�^��`E�2�|�CVU��6d�M�����y���B���[�ؚ�&e^�l&���d����l�EΌ�3H������������$��۲�S���,LWi�L;>��G���Y��R��5C>.�C��ǪAx�d4��A*�lL�a���f��0��c�7p��	�M;Y]�˱lr�A���d����K�F�<&��c��Jad\0�Xv��4G��aN�sP=�$��]�r�;r_�y��33]���O��=�6p3��AE����I�D���� �]��~^�n���CI3,y�3����}E"�m�
OV�W�@&,��B�fw��u��GY/��L��f���e�4���$2mM[D/���M��"pu%i��ф�e%�ڶA�ϋ`ZW~K9�����rO\�f�L� �Y�D�;I���]y��͡�,��Z�� ?�N#�nE�i徂c��᪞3f�jː�5�Ad�*���hG���j-q�#� M����K��ts���*9�T9	@�*JM�4P���@�2�',�c�Z�t2���S��պ��X��̢rʉ��`�]$ɘC�`F��#N��{Qw����0����WHv@4��C���V�`�YY�Y��a�pH�-�V�;��TI�6hE����Yu�^\�6��۱� ��-98��>��Rx��q���V�B�����*:�]�$$g��%�8<��'Vҡ'�k�[QE�*����B�C�S���m�!Ȭ�Mh� �p$'�o]�7j�[��c4^��4Y��I��h:����L���#O�]��BACl
t