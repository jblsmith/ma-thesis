BZh91AY&SY�u� ~_�Py����߰����Ps��]��u�:�H��&(���FOMC!�L� i��I�mG�  �  42&�*P4~����f��4@=@ 8ɓ&# &L �# C �!L$dɣM���h4 4 ѵ$�i �B$�B��!��G�w^L�4�hRk� 2Mv������`0K��`$��{�4��Ǽw��-�]��4Ԏ(mzzp������idd�r8}K��إ�rJ,df9#Ɍ��O�i�$Y
D,/�M�y��9qm�*�0�5T	�Вůdء�9����}�F{l 3&M��ؤ��G<,�A�H���	A�Z��3��5X��^�LAd\�U;�$ȿL_�,�
��� ��c+*3BBB1z����H���3���jЇ~�.�N`���h��xŚ"/\R��Z^���J���C^��/�H�U�ѩ&t@�%$E�AV�^�Fv�62@M��uUG�T���p8�Ay�M����m�@!+���v�D��XP�`�w����1b�6�p� �?��E-���*bj�1Е�*jMSjÄ�A��w3��K�h<��t�,)�[<�Kz�y�dn�K��N"�E�,��w���.0�Z���2NN�.�JQc�����}��\�n����~�33 ��	�w(��cg���v��-���,���C{�cX�b��@(�L ��i-22�`� 6՜��q_U�DB�dܹ������WʼC��5���MN�@p��\�r��c��2\�i��k9��h�����@�5`Ĉ�?�(�1ӕ{�q"6a�V����v3�炭�4�@49���ZT%�qQ�xP$����#�ref0	z�{̠v�L�)y� Yslc�������iM���㍂F��l6��KQg3�&�F���b�$�MO M;�P�V�[�*�M,�*�� �3���0�u��\����$�G9D��0|~���e�n���d0D�^��wE[��V���z�[�>S�H�lYZyNc����� �g��HZ�&�rH7�l��C��#	�R����QKh�;�!HJ�HTIըʌ,���9KOY^���bҦFp�A�񾖥 J���n�\��r���Rs'��0���!Ƥ{aB�����0�89wxob�n	�7�:�g{2��{2��~�f����o�]��BC�m��