BZh91AY&SY�ϸ% +߀Py����߰����`�dh 	Hҍ6E=&��� � ����4�MQ��ڌ���&���L� q�&LF& L�&@F ���2b10d�2 h�00dɓ��&	�F�!�*H�512T���E?�H����<��P�z���^@��$����Dg'�TAy
��'��*}�&U%�+���K�0��c�Y-o�&1$�I��L�)R{(�K�ٿA�n���_w**�~-�g�ձ9�s��'�:��!���L��+&,�C�j�*��0
*
s�^tC�!)�?)�������K�����R��R��"a;�H��x�<	?Q�n���m����nӐ��� v�9����²��0��D�=��ާ�?	�/����d����c�=o��˩���UEJ˱���fS�U���ܝ�SmN^o]u�K��S��ꚜ��L��ȸ���6�<7�MŪ�]�E!�Æ��Ad�� �Rn�G��k���tt����·#=��& �
��rNRu�/��	���GE�29y�x$�(�'����o1b�n�i���D�]�h���AuDV9�q�z�Ƀ%�7$��6K��R���ʑ�l��a>�`���srSa��0�Y�ű�#V���2��w4%�hy*����̏D�B�uLYEw�hMa�7g'q�%���:�x�<bB��$�C&ffq��y�4�i�����`�4�ং*~w��2�q�_��e%?7��i-S��eU�eN�&��K�1T(�i%�F�)2Qz��u<
uOuZ�+���V_��=4��j� ��i�9���-ba<��Q ����2��v=�����=G�L\j0i��ϒ�(2�������#=�I>g콇�5?	�[��֊T*��E��h��d��m��Nn(�L�j)y��d���\y}��#�9��$��/BD��ΐ��"ٽ�l��'�����Q��1?��Yg�h�%�2��n�~�����g�;�/RїN����(N2��T���xQS�(��f��k:&#�Ē���۹S3&��'�3QOs�M�:f�M=S7d�(��s���z�|�nf���Qb�I���c�Ձ�.��.��\��d�_��e.�*)��䞮�{C�ńfu��#���8��ѫv\:Y6�bI�j�R��ԥ�}���Ɏ<��CCr�[��+H�Q$�e��V'�OүU��M��,�ڲ����2c�t�3F
a/�t�����Ϧe#�0���&�K4,R�O�Ǚ�N�l0gVb�v��.�k�dy�X�Q����䒻�M��sb<�LX�C���tБ�d�Ph������c�;J`z'�6ʑ�J�&�gk̇������%�Ǜ&�Y�jorqhj��F��J�,����1`�ט_I�`����;W���5*mv��0M|�F�l4���S<Y��㭨g:3��cL���/ƪS��Ԏ�K&�N��um��֛Z�ݫu�m�%����1��#��`մ��89{<w*t7�N�GT��c�ݺ�q�e�;ޗ�d�j�'$4�C�]��BBg>��