BZh91AY&SY��-B �߀Py����߰����P�q�'n6�];H�����T��j���<���=M�i��4đ�4�@�A�   %4"'�MOI�L��=@�h0`��`ѐ��&��D�ГЏI�i�@��@ bi!#!�F�H@��	���H�b�@u�u�����V�@X�9�t�rl^���ko���ϑMQW�߆���!�I��
������v��\���=���������wb|J�H��C��V�@04��������Xgs�p�f���8>��3&M���F�_��;�5c�3�W2��ZE)�ID�K�&�X���d�A��sZ��ұT!ځ(�.2T��VO$��{
fi%Z�]��f&��b�B����@�Jb�"@��䴝\�\�4�)e�m7����[�p�rSǫ�1�iI		.	$�3�O]ۚ;���1$Tz�y��[j��MKm��p����* cY���e��u�X0(d�S�V�@���wt�&Gl!ڵ�b��y�{����`�vq�~[��ƢH�3><ڱ�i�l����55���G�# �$s<�=q�>�ު�W,���}��T3;���p����F�ڑ�D�S�~0�QE7����K��AЎ�}�4K̬`[2P�<X�D��!^�\�&8 �D�R��xL;6Z�e�C�b�/�&3j���t����^�8ˌ�>�4�K*�ڕ3�s�x,��U��s-�Q�銀b	̅�I^�]�+��;�dg�Z�$���TG.���Zn�ʚ�fzs51�L����c{��;1T���6� 06���AMfѱ;6��kd&����5T�h!RX�jy�h��%BBI���ݔ���,`�B�8��G��M21����.�Q,�U�5M��{x�z�01� ����%*����)�:h<��8����.l`֭ds��L�1Vlb�ӫ��2N��H�--N��~+Q��v�(�^(#V]�t�����7���/�e��.�k��4db\��6�(�8,m�KD ���Md�N�$j�,�]���\,���tR|cA �(Z>S5K���ջL����/u��2�e���M\��L��zk��.�p�!��Z�