BZh91AY&SYo� _�pyg����߰����`	?}X㎰ �q��JUR�5O&�=�F�� z@ @ڏP� 	) P   4  ᦙ�&�`L#��i������F�  hd   (�ME=��O	�OԞ�� �j ��Q�x����=2z"i�4��z��� ɣԨ
���E���!��2G��EnA���~#���-�@�0p�|�HV��DH�ɭ�a 8�Q ��;bT+Ah��%�f��o8���Y21��d�Q"�7cM��������"]�F�	���Wab�ע!�%&y�ZH+������L�l��N��m��'
*�#ɬ��y<�1E��z��u�#��w��nu��^i�l�[%��i����)0$U����v����Ƽ��mH�K,Lc�{<!7�����D��a���+�璁�қM̲���b��TV��E �J�g�#I�$�	9㧨��A����V�xkz�n���5M��_��u�O=�υ0r �,gU�����d�K����tp�գ`�쐴kz�Elի�$�P})FN1f��(�6���d�u��UWS�Y�.Z��	�x�	�$��J�XO�s�XXB�<*{2�Gq�!�r�΍xt��j�\:��4 ���f@0a30�jԵQS�.z(c!�t�� 3if�9	;_%ZCk���,0��E�HJ�H�P�PD�X�V�1�`�Aѡ]��:�K	i~�}%n�n(�	%8D ���=,�ࢣ�N9w�E�����Z&��(:B�l�O��f�����w�᥌�	kهy%�@4�Gp� Q۪29�|/�W��0� YA�Ю`�C��z<�����{�v\�a�2P�nR�$����B�����
�]3��1�M�껐��XU���-:�v���pU�
J�U'o�������à  A
$�{0w��.�HT(ܱ4�5�tJlة�ʺ�J�([�U�%JRL$�� p� ��@���������b!�'' �BQB141,j�)���H�J-ik�cWs��ܛ������&l��z�/�.��t� ����M扱�[k��A��Q�:E��� (Z�G����@춊#V,��!�����6r�r����x;��nj_�[�v��{��Z�*� ,�H�J���`�:���Y����P�BQ�X�B�?�����C_;L#{<o�z��BOo1'��������
0�@�g�ٚ\�N�а h��$�7F��@&-� �Cu�*�ho�'nԴҗ�n�� $nJ����m�ѫ �
7�@�W������1��=FC�Y ���U�T	LO+�N>�!���F�:�'=ư�GJ��;��-� ܿ.��=�/���j6�9<��
 [�XD�Ibs�\��'�^�;9㺵]_3�Q�w�?9�5�r�xzGq��t;�@�q3a�Iף=Baͱ��v .ǉsa���a�O�Ɩ#�d�bs�ɠ�P�@�*'a�P8|�yi	Q5�G�(��%�6�C�l�v�����E �t�+ߘ`/�U�	�XQ%���R�kD�7@��Ҧ-�
�5h�(5n�aj2`�Qh����:=�ܢ�A��8<�y�Ft8�k���a�����������^D�02�P�;�	ܺ��=��:���� ��w�J�HՉN�2��e|u+w%%MK��ζ�r`�.	�*\� ,$��o��5}��ь���<�6��&��W��Ǖ�x3q���o��������Vq��a����!Ct@C�����J���f8�] q8��'aL�Й%J�Q��ܭ�h^7�P�$�	�<�?Xn�@�f��ҝ�1C��Gc[�x��
u>���^g?]�����ܑN$��B�