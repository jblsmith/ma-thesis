BZh91AY&SYq� �_�Py����߰����  `�1 �i*�  A�zOTш@ �C&� �L�H�M2i�=Mh���4  ᦙ�&�`L#��i���$��Q�4���2 dh Ѡ�  i���i��4�0LL�� �" OH�=CF�i0# i���7�BosH�)��A�Y?���Z�N?��_)�W�kk=��Ϯ�أ�����3��.�¦��Y-mX"M�2T�H� �$�@,V�5r�Dp��&fi��B˙��W���,���\cW�{�e���:Ohٱ���ZTR��V8�,G#wʵ/6g.^j���I:��[xm�tNn
�E0s�2�[/+�
]�~-���e��y�g�D�璮Bm=�s5�?\}������C��g�E�.�k�����(�U*��e��fS�U�k����P�T�k֫؁�)S�)�U��#pQ6ݣ4�
�b�B��T��$�ȸ���4Y�wFe����̜&,Z30�I���F`���%J��h'6GeI�iIo��TaK���^�Q�d�$�KC ���I��,���NS2	�\��똑a��(���s%e�0�1$c!�V�Ud�y\��L�MYdf*$0�����Ѧ���x��Lj�6Ζ��0��61���m��!�ɛ�A#��l�#�Xg�C�*@�R�<�%K݂�L� klh����&��RL���B�mS�}4��*(�b�ű�u�j�uWf�0]��b�s�.w̉ի��I�@s����b�?	�<�.�K�A����%̶��k��ytӓ��oË�����wlm)i�[^v���~�+�kg~��Չ��mR�[��F ��;�g2���RP!�=L`B3���|�>i�x�~3�N݈�2��K���N�@�UMρ�B-�\���L�(SmH�y��%8Lf�<rě4vO7�|f��ıe��i�o��{UL�2��v���'j���t��K�Z9_U|]?U�)DƎ�P�����a7Q��Y�1�-��H�䊶��jt����Զ���h��S��Me��9MZ1q�*f�Ƭ7�z���/E��\��X�F
`��j�䋳sˬ��lvw4��{Nr�W��h���}���'ń�so2v������S����n�o-�Y#Y�J�Eph��?n�z�Y�^/�yG	�"K�=l|ޱ<��U�^�$�)s�Y��e���2c���q�ļI(iKw	����ua9���)K�\�����L�e#q�uf-�Fic�vk^�3�1	c^S��yQ��<\N/��w�=-���E��͏)��f�m����mq,7kgs���*��*&Ϡ�硃uH͂�5�v1�y��!IF
�)�f<ċG��͜�-�mj�w�M#���q�3T�p��9�:f,��a1�I�`�S�s;����4T��g��0M|�#��'v�o3\uh3/6��[}2$b�qp/�U)�����
.�9K�㣇Ʃ�Ͻ��uKuh�7�%�I�e�m��v���:W���c,j�M��2ԑ��-�p�Ym\X���(6O��KJ �
ЯkK�]��BA�?�X