BZh91AY&SY�
�2 �߀Py����߰����P~]���*v�̈́�&Bdjz����DmM�� 4�H�i��j424   �   bi	<��!����jh�M  2�L�1�2`� 4a�5�i�SL�HhA�@�� �q,hE !*���'��	��V��L��OĸԉFkG��deCa���/�x4�C��~$ ����^���Tp6�*�7�_�o��Ab��
�
<o%�H�����/����̡ֈ �Ƃzݵ�u��'�j���ݏ��	�2i[,X)�lhZoF�CR5��썁���&����G�@J?���n*,ؗ{�j�L�	F�8{�c�$1�jȶWt.-�XXڋ��΃x���M3��W�A����?_X>a�I�KΒHA�x��_#��Hu
/�w�[��B�,����?���!@PXl�$U#�^��@U�;�=B	9�5�olzr��ekƸ`t�1U9ql��˯�h��aA(��"��_/����*^7~L�_��w/���%JCT\%�W{�ι�nӍ�Q��33$x��'^[E�c66}�[�(�ʨQ%��J?d�������Ώ����n$��ʁM 0�SV�uV2����ߪ�T̞�I��h���p*�!��3��t��F;m)�M59h^�F�*/./%���!Sn�T��%!�;r�h�d'%NM�uAu��nr6��p`SL:� �)��+�����y�N��'��-����!Si�fR�ߞ�:,��
�ͱ�>G߻TF�u�%
�
��8Am5�
�KIO#k�R�E���(�%N��@�)a@
�V�}�KMh;�!����X�8�f�(,�r`:�F�h�&��sp�.����"�a���S�l��!�
��4⫥��l;+K@�!�o�f*�+�,�ƅ�L��T��N�E���9�~Z�J�V���!9��&��	�Ej����k�7�Y����%]�!�b0Xme�DR�
Ec�f &T�J��,��	jSM!��;�$��1:	E" J�X�ӧn��Wv@��i��׷=���4���k���h4�բ����)��W��