BZh91AY&SY�5�u 
߀py����߰����`?k���y��@"���Q0S�6��4��@�F@2hh  �	�*�` �0  �M0F`��!�	�4ѣ4ɑ� �HST���h  �   H�hF541)�4���e  i��!4)�4��2i�� 4�&4����lAB�WT=�F�e���� 
8�c �Hs�ġ�����
� �Ѐ�i�� �d; 1�6��R��W,�����������(��S��K���pws�W_���5��EE��BꄡC@`�z���v�{Q��!(݃zh�ɓِ��`b�ݍ��x����$A7�L�EK$���N��arOt���_R��9K�R��V�����3]��v$)���+�2��l�XI��p,�c���ׅi��K�X*��d��Η�;Cܾ�<�^s��\V�{|�}g��r��*�YN�m}i��'��Fgt��lD�/9�L�پ�3x3	U�3��1��WT���j~�^.��V�!M���7��(��G8QrP|h�Jl��XF]4j�mF!�.�5w�X�;�P��[#$����ǰ,���.�f�i@�*�NT���˼���Z�0�V��� �<f�֌.�
0�u5���/v��b��eP��4�1
Y�.�9�1@b� �Rhj"��1YqAh�呢(Nc�AR�Jl��,���ك�(���Z�.`
8
^�XfN�VM������1�.��̛l���%ɘs�;XcŨ�ow�
���̍̚��(�ʢa�牧)�w��*4T�f5�(����v�/�x �t�HFN��I$ a���R�k^.������gr��hH�����TiMʱ!m(��"��!�c�FD�&H������B�rb)(�'k��V����9��N6\ϖH��#�l���q,b��@t�S4�9�/f.fr�S��R�(�JMm�m�ۣ̍h����2��ӡ�I���~uc�����"v3&��T ,ª3���pJ1�~�b7���S�H!�$����C���z^�XjW�ɵC�����)�,rr���,���o�2��B�̇��Q��N��9.Y��;N���|s�H$�mvd�=ɓ����	`ֲo���9=�w1X�FlM��iN�C��gw��n@(}�A��V�tc��v��zv���AAT�`Z<��F��\Q���߬ !��otr��r[�SM/��h_�`��xWk �T��sC��'8�pY�<k�|B���*Kg�zI.yTӱ�/fM�h������If�M�Z8��T���1���{��D�-)�(a�H9�M�@q�%Q�U<{��&,�7�v��8K���`�	52$�����
��j���9��pGz�,l)~]�_Y���n�NѤ�$��s@�6���96b5�҆�ڸ���i,���ÜB:;��*����4�6v�M�b��JT���JP'B���J�i3$n#���Ǩ8�8����
��;Zd��pH�o���U$�{Z��Zfn9]�N	�zlmL'��` 3	"L�v�PQ�fN�6@{�a�ϓr^�gvݏ�X��~q�4z�mN�����j�2�
������I�Qj��	!��*��Ž�������-�7!$i�h�5aB��e���`M�G���㥀Ş�2�j�d�[��CM��67�o[�3P��º��=�=��.�p�!�k��