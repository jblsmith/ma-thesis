BZh91AY&SYO5Q �߀px����߰����P����E�A@E0�Ҟ!�M(~�Q�����z�h�"�!�� 4 A�"i �� Ѡ  =CC�0L@0	�h�h`ba�HhѠѣA�4 �   )$k:��(@@ �	B����У��v4-�%���ꐖc �2��89�ݲ��O!畗7� ����O�A�;����H���\U6�VE[������ ��jy�Kl[�`��
�A+����>$�!�%`A1�� ��@Ee���)�!B�#*J��$݌�v��\/3b���|b�Qm�,�{�hҫ�J�����U�� M6V�Ԝ;!+��Fwׅ�U�qj^�V]q�x�����&	f���
F)dց�"�1$D�Jle!@l�� �F��'(=�n�U\���<��q�֟��C��66���� �{��)�g�(��E9{�+��$5�L�B7��xl�=S oe��A1l蜘]�j�ճ�@����]]��(�)F��
�]�rؚ�����U������{�?m�q�5��~�Kn�{Oշ���Pؓs:�<�[&kMI�̵~�O����lC2A���	ן�^���_R"��9,�Ad5n��Ki��H=���9�����dT�v�H����*�X�^�Y���U�=���|�s��`�*���̎J��f.��L��i��ML�ͮ�QȰ���H�.�g�	�?�0ǎ�,j%]0&�)*�P�V�G���trN�B�N�+US�,��2���BtV��wa�Y��f�Fc[Rq��r�<Ui�4�0�_[U���JR�]�S�i80�� ����.����STM�:$1p��R� �@�&Ĥ��B�}�K�%�yC���l}lH���Ōd�*	ĵs�D*��ۘ��ۤ�RA�D\/.EUO����+�V0��t�����W3���*�LE�! $�[�Be֜�:�@ߚ@�9V4�tm��V���� �	ʪ�Ձ*!TUMC۴�VnZ�d���U�_qaB�4�3�4L$[.���H'h�T(�0��4�M_u�Xk����AMtR^� �"��o� Wz�.�콋r�`��ۭ׿m��	c��g?��bɐco���w$S�	��U