BZh91AY&SYyW�W r߀Py����߰����`��@�a� �(JyS�H�6���i��� �P�F�Tz�@@h     �����l� � i��  q�&LF& L�&@F ���2b10d�2 h�00	B4�&�d��&�h��M5% Z����4
P$$���R�8_���B�K� Y�X&0m}P�ԹL�����+T$6%�bƘ��CBAB��Rb��]�/����Ϣ����s;K�!�
���2�C9�g��z�H{��J$�8���3�Kh���d��aD �M!�u�E�� S�j�t�=V�B�rM��!`���̈́���/�_�����	V�"P�f��|�<_{�,S�^�G���1��4$6��+��[�2�AQ����`x���{�d���T��|*�y��d�X�x�Ah,����g�]��cP3P�{f��(�X�� s2E�+�Ow�lT�-6~j6Qay0�CDd���H��$Ł8Q\��Y�DP|�h�$�+A*I%B"������r>]5;b�"�F�R�l�E�+���(��%���h$�R�N��uP��o�N��������[m�&�DT�`zBO|�i����H���Xj�m�`��^���6��3�-.]a�&0�iP���%Q� !)��	1�0��z�p�Z��p�]�\P�E�yT��d;B�����0��K����~��tf+����f�O(?-�S�Х�2)�q��|��2D���M��xD""AGʾ�q�#��B]F"Б�!1����7-�נ���B�*��@>��'?�g*�:��w��$|�,�R~��8T���4RAcb�W�f�{5%	���\=�B8K T�r�)"�'�f
���4cx��P����8�Pc���Ă�P0j���a쪃�2�h�2J�#��!�EËp�����q�47�q���\�Ȳ6�X
�ĝ~�tI����E�P	(@vC�؉.tې=�[��`�wx��)�t����2���n? �t5���z�aS@���MCL�����
��V���7��l6.������;� 5����>�aD�!�T� `q�����Y4������"I01d#�Y#�Q�U�L�  ��@y
�m�R�
�$�"���,����@P���s	>9�n9��T�a��s������r�>3��dh~�;���M�ڎ1��A�*�04ihHȃy^H��PpK��r�"��,b���3��d#��c:Q�� ߰ڪPW�I�dPvZ/�7���0`5���eAc�QuKXj�/R�AL�e��HѕBE���E;�L�m6��5�kb�6顉���Nq�i�P��"�����=ė�=��Lm����� �2R��+�]U(KP�bٌ� Kp��q���ٝ����)�ʼҸ