BZh91AY&SY�w� ߀Py����߰����P�#wgLfݸ$�LT�E?"56���z��ȞPѦ�0A������&h�i�  ����OML�OL�h2ae?T�2dɈ��	�����$�2i44�4��    =L�	Y�$�A�O�����f+4�!����N��� �G��h.�/�Y����7�9ߎ�%�"���I���*xϕkx]C�<��oG_��LYf�F���dV�RX�C�s��0H�F}&k��8*w�-Ze	,��d9:��7i���鍹Hm4��ſx9�c4=�!zY����8�9�
*	�E�J�<��b�2 ̋��^�T�@��H!��dX�b	`#�:���[ d���1k=��U9@ΰl�����,�nb��础���V�� �구�n�a��%��EM�����;����66��m�IA]8mS��::�&刜����u3�Y�����t6۟lX�����^���V�Y�]��K�C(�
��-�s��~����1Y�Dt�k������]�'�f��$��ONlS�{�T1�U5����}�����.�mҔ��*���2����tc��a#�p�'/��k7��&r���"D��"{\��#�}y>� %o �ʍ��le���
�Y yP�m� !�N@�q\h��K]��MA��c�.%�@E�>��i����1	��&���dΦ�$8�'(�x��+���)A�)�����D��0RH��'%�Y�Q���g?p0�,��$Ju�J���}jC_��ȑ<G=���0ǜe�$L��i�^���X�=�fjb�h}Ԟ6��i����f�� �#p�i�+�K1W�-Pd<��78v��+��Ҩ�
D�x�$@0Ő���)(-Ą�3���B�V,a)�(&�-\�B�kAƿ�W�k��}�Ch$%dO�y�И:iH㞤�Q�q�����̬dtM����a"d�WfT-Č��`��k�@�b���S!�sܳhE�̑k��*��ɒE�='��pN�U�b������VF �H�Y�3��*k_��"�5��P_E��b�~�b�4lY�r(dPm�=H��_�����0�j���ʃ�Y}�]V�̰���d�j���L����rE8P��w�