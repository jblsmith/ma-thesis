BZh91AY&SY�e�� �߀py'����߰����`����1��  �sL��Lф�hшd�� A(!�I@f���F@�@�z�4�5S'�J�#@ �@b  $��54� ��b  �220CFi�F i�# ��#Bi�D����Sdj=OSІ���Ꞛ�آJw��%B]$E�CT��D��i�M����U>v�:����4�"\�¬��j�k|� l����*O��TB��LY��J��'�IAO0:u� �a�)T��Vq���9bG��Ë|e�mP�BGp�L��(�tR�ɸ�n��n9��"rg^R�H!�{���Y)oߒ�޷%i���&m��^jZ6y՗��N�/���~m_q7�w�$�-n��d.+���Xa����^`�N#d&D����=�Yk��*�lvۺm�����d��Zb�d�aQ��w�¬��i٩��H�͂�J��'9D��X��Ij%CB�$�̎*�h�!$��JF!�c*NɊ=�I��yw��1D��'t��H�$X��E������PvI"�,����L�"E�ČՊJ����+��3����J�Ñ.���X���'
�\k��FJ���R%ellz�t����F$����OE��� �.3�I<sc���7�=��1����lLHPAIzgH�!Z,*�� �jCܙ"T��&R�
r��TI����/��58���B��H��a�/#�K��QE�D��h��Z�%�It-;`�J�/�vG��0N��u�y�l� 9C�d>�6χG������G)�4�&�k��7k��k1���ȩ4c�k?;&��ƾr��c#-�\�'�9~t=��R����듹�)DO�Ҕ-o�G�sO*ǹ��ޏ��&����,�8�9����Q���dO��-Rӓ���L���������0��ye]C߶�Y�ll�2��m��N/�GԪp5pƗeRѾ����g��!�L�H�~�QSk͔~�w�����0�ԉV����S3'B�gz3QO���D�M�S&��&i�r��o�\v�'�cf<�D�K����M�H�7n\OS5��r��0_��������䞮�[C�Ʉfq{�����p-+f�l�od�t�4nR�Q\�J_����^�8�yJ�k7-�wcdAۗ��7-#���W���M��Y��e��ɻ(���S|�E�
�h�o�H�D�y����S�X�c�՘�]�-�勲Z�a�������v���Sq�ȉ��x7��u�x�O�ۓ��g�d��n,6{��tz��P����zY��uJ"j�t���x]V;���%���d�+6�Nwk�CTu�7*kYg^�\łu�a}s(�[���u/ϱ�jT���w�0�rHm6B�3%"d"ӱP!1�h��&n-�i~�R�[���T�nT�2�}ۚ��k������ͮKCt��șp�Rg-o��缡���SG��h�=6>�;��)�_á����$ਢv6}��w$S�	�]]�