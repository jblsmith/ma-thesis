BZh91AY&SY7
�R �_�py����߰����P^��p�ɭ�NIOF�	��I��z�MM��z�0�������4��y4	���  @  ����SMF��L�h��d� 4 � 8ɓM0�14`� Ѧ D�De3Jy�y��SA��z���  -���Ad"Bt��	Л�t���
��I���^�umT��"�6���ʣG�����F|^<�ۇ�3?n
-8�:�EG��vۭTj���We�Uօ8�F^��M��%L���
��������ה��4�\/�B�[�C��C�o�����a&dɤ�N�p�؝���Y�8l����AP\ki"�rXҨ���`�1daF�3"d�frE&��@J�rԥ��u��GDUYJ#i r�C!�:�D�!�T�,4I�z�:%�G���\^,zFI�[J�������w�ccoe��4�S��jye]	d����Z,L3\�6���,�Z@�Z�
]p�7���j�g�bݐb���MdО}��lp����]���J=�m�
	���vhEn��;i�b��p��^!�O����ԗ�[�b�����K�fBf�9�N\v��Tjl����G	R�5∹=Gۛ�c(�Q��J�ih�	�J��)�%�Y)��\��G7(+������miӜm[Id\�v��Hh6�J	�MU\���Do,2�0&zɘhbd��R����x�\���y5B>L�r9�Uzpa'�r�/,���.5.;S�:�����D�<ز�x_,�%2�`h�F	1�%DD��S35wۛ�x�'s
.���6�p�gtV���on�T�h<M@�+�"9"��"�� !0���T�D���'	�an�afT����hTBOR8 t���q��!��2Z�Ģjʑz�4<?�pCAȠ;j�Mi«��6D۔l<+CAy��d�,bW���L�PK�� �P��xБ\�m�+SD�ʔXb�8�]�S�I>�J��E�^�L�
ߍ��Y<�
.��#]Zf#ϖֈ���5�"�db�J�)@ͦt�?~�����̆Z�.\F5�)����H]s���Y�$�w������:2���?��H�
�]�@