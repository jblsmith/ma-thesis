BZh91AY&SY�I � �_�py����߰����`_0�   hh�4i�F�&�@   � J D��6���& =  2d�L&F@��M#4i�2d�L&F@��M#4i�2d�L&F@��M#4i���@�*y6�ا��3L��hhd�3S��Ho�d#5B]%�MR~���0����p�����J���Ҥ/*O��K��Q�~�Ւ�у��)5JT��@�0;����k�9��&��&�u�}֛�����s8:�XX�9��ַ����W�Ǐ����|�\B|~ړ��\TR��'O-D��#^EeσQ�u����b�Vu���V�c�K��m�U�V�V[u\�͵�)��RѲ�e�p�f��5�/�O���kK���� MS�~�?U~'����˕�I����?��m���*��a���gٮ���Z�7[�m��N娯.�擨rD�FJ�=�xo����D�2Zw���(��Q?�����k�-;��n�SҮ�,d�J���$:�J�W�W������	f`j�k!��7����5J�s��w�A��}��	�˖��5O��qGETc#i�5
9q(R�1ud�sq2`�j�W"�Q�m�6�+��wc��0ٳO��ԫ$g#y������T2���2����֯ӭ�T+@�`��EEcH52�lX��=9�1 ��Ē;�X�2�]�J)%���ti��G���q�٫n9l�fM�E�:=���~�R�JUsUUURR!e�=����ۧ�����Y����h����԰�������I�0T)�-�%�Z���+Rв�в�����ኢQb��-l�Rd��1xM��(��O]�گ���2�i��Ǝ�*��<��d��lp��?�O#���7$�h���u���|�pl�������1�q�S��b\�3;8��^�O���7��#���ϸ���~��I�֊P�괥G�{dx��|𬻞��'.����LD�����uD��iJ�O�C�;T��K8��N
i%�L�t;=z�͇�dK�(��U,�G��5�K`�+5lg�:^mx�������U�ԴaɆ�t��]����TC*H��l(����=���Y�lw��#�B����Ω���n��E<\Z�)�fɩ��f�Ƌ�TyV�򱋕�ǚX��L_k�Uby���t6k�=E���40�UUU����n�2O����ja��q��)�N�Ҷoǣ��q�!��J�Eoh����)���q�;�:���F��ԲDP���<�v5y��I�K������ʼ���.W)�.�$�E�"��Z>��)����R���I�0u�z�]3�X����3�f{I
����~D���7��K�������>�̞��sSqa��g~=r�y�D��w��q2]R�)��űC����v�3�B�ߣ&�Y�4g��t�i��n*T�,�ξG	��y��t��GJ�5��6�s��&�#��k�͹S<Y��4f2�2�-���f�r7K����ppGK&�NI�g��������R��7�%���$ǀ�o��>�Җ"�/��	��II���e����Z�P�H��QD�m���?�.�p�!ƒA