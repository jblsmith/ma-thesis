BZh91AY&SYY�� �߀py����߰����P>wWZ�0v���tH�hL�Jd��f�i4��i4���@�i�Rg���@ �#F�@�2hi�����4  sL��Lф�hшd�� A"@�ii6F�4M4 �44�`j@��"HBPW#��GУ���ys��+�HbՒ�k�vM�a��#d`1�wڍMh��N�_�DN|O�?��ꪫ�O�i2�i^����f&��7-���<�e��,�e�N�-?�ĳZQrP8�4*�HV�?�D��D@��T��a��uN�1g-o����� �&���w�x	$��Ro�r/�[�����t����_�
3����[Q4���N��Y�&��_ݗέ�J �]\��=���XS��:�L,j�*2�j�6m�ƞw�EwNhL���O���8���j�C�=Ճ<@�l��)�θ�`v<wcv�tT��l��oQ8��f�h�ܐ���N[GR�3:K�c����O��r�Ff~��`�!n�]�^Gw�X�%j��2σ
��q�Q��P�10��
t"�%R��V�0�5}f��H+n�)n���4uF�=����rKw�Ǭ�\?�����k��J��L�[C��Q�x�����EVX�w�.,^��3F�~�M4��2�嗲^U��y;R8'F�9 <�$�Ŭ^ⳍ�q-G��QL�NR#�I�G��a.��>��	������˘��8
h8�t�6Z�9!�BѼYus��60W�F�bi��4��mm�,��Q�6�7�ܜv�E����4ז��cgS9�#��`M��H�4�2�w�V͛��1�,V���*+�d:2����\���i9$�\
v�\��ȥ��:r5��Dqݘ��� D����1��vD�\v³"@OS35�3���P�×֛-u����$��è�,%�ű�I��㑬!P�C�$Rjy�h��J(4�Y����d��aP�"q3�-���¶N\ʓ�(%X�U:
!)���s���p3�1Ak�+C�L�篰���:iP����S��&9�`�,-�&Î���э 1��<H\I�p��5iH\��u/���ݽ\�5W�E�B�4e�N ��AH�2�mT�S�8*� �� [Q���V�"g�h��2�umt�5#cM%��Z�Xr���y� �Tcx&����K��*.��(��я���0oT��ܺ�V̱�%݆s�[�\ɐ_����c�rE8P�Y��