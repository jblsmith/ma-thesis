BZh91AY&SYiK �_�px����߰����P�s�w�S���V�I0��G���&���S��z�C�d ��4��LPi��� h �  ��I�4��F�m@  �2dɈ��	�����$H�&��T�=LȞD ��h�44�H��@�Љ! ��%�$(�$|9���P��"L]�A&���TЕ� ���c8�Lk&E�.זo�y�N$z]��xچ��N\��������T���Q��X�X���� �VA[xЩ�$6b��u�v Xc�d�K��G���+x��\룧�]�zj�ǩ�юQ�by����c廯��M�-}^��A*�HPR
��t�\��%o��a���.,���&�f�S�IU��/Zwy,m�=y-[;p����jh��dY4��gZ5��1v�^�z��ԕ�8�+"�Xw�� xU�er��(�t+�nuQM�d���*Ğ-f|js-  : ��:u�G$2ǲ��� ��aQJq��~P't K�V�K�i�	.ABJ�5
%d�+Q�5W�����o�{��Y$���En�[�}s8��W�����I��%�.�ME��/��]n��P���}}�d�n�Td����5o�8�doy��#\�fH?na�r��ֿiftM*'�!]Pƺ̊���w��#�jAʎ{ ��f&wZ% m��k�W?E�$CZY�r��ټ9Z�9�r�9�8֖��`ң�yu�40��ZF d�D�S�FFzY��r6�ɰ>��J*�ز�W���1��rh�+)n�(��HQ�ir;\F�����A�2�=^�&�b�n:UD��tPG}E�s�f1CP����� �335,�s��DnH��U��ؒ�$��1_	l-�=�jah�k��Cp�*��`� yITI$�X��K�)X���E$<��s�ީ�ˉ���ʲ�L�'��e!�!7�K�5�PY� �DZ���ڡ	vD<yry�C��Jp�Yy�[��x����g��m�+scH�ꅱ�2.f�@d�E�z�l�U9��IE.#�F�$rH�ʹ����*�6Sr��4๠�֒�ޝ���ጮ����#Jx���!\̥Bek�+Oit}v3����@㞿�i��Z��0�j�ٲ�3h�9�M�[�2�C'e�w9-4.��w�]��B@Tm�,