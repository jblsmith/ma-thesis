BZh91AY&SY��� �߀Pyg���������P~9�@�Ɉ� E0Sjf�iG�z����f�T=@41��T�A2*�4 4     �a&�BSM=L�zG�4�M<��h ���L�1M00&�#��M A"I������z���y2������e�	��D�$�J�s� I!?��:8 ����s	"��@����7����h&ҵ����4k��8������I]�����������N�1�c��_k[�A�ŻM
�^k� ��f��>Y�ͮ`Z�e���d-8�n�A��j!����]'*% �Uy\K��Aj�N�$��MI$���C�ؼNGa*~<YYq��<�F��!�2ho�<UpO������_'�wxn}��:��WԚ��(���$�gY�t�o�j�M`Z���3e4��(�Or�=E�[˦�k33*�PQ�p��U�jGXkb�����Ͱy`��ȹ$�&�Y��m�R�Y�^R�D����DF,0��AȪk!Sv$>W/ �"��J礼����[�qy�t(�f��W�-��%]�Ql`>(5�a\"��k���H��s�gg9��H$YRI �0�9n٨�����(\VG2�Qd�C CA�:&�h��	
���"	�!��e�a�dQ�g�n. ��{zص�y?*O��믵��ׂ��~�������s~^�m�=��w�M���??m/�k�Μvצ?(�nz����~.��B?%���.��F��s��D+C2|fI��􋸸�o��ׂ=�ȥ4�+���C^�1�	}�M���T�#�AA���T��"P�wƍS�Wm�K6so��n�of �^J��1��u��i[�)�[�4�z��� �ID �mMYY,L�č�Lg�p ��Y�iL�kJ�����yKJW.r�5q,�mi�~.G�Ї@�t��%I�,�'�Z��j�D}=�R*G�ǘ�F;J�MP	��6�g�>J��kaĦX�bY�36�5W��(�lc�[7RcmkۚA��T$W G{q�Y`ev��j�Tr6)���I�5;�h��%BHBas!y��b\2(�:���T���,j��\����b*#Q�$�C4tzy3�����u�N�UT����'�V�W	��os�h�ꍆ���g��m�6G���##5�q�I��@ՂB�á[K��uW#5zH�V'm���m��U�(5��*��5F.�wr �n�ciYyl�q��)0�d�stI)h�&�������X[l�9SF��(]D:4���X��e��Q:.�_��,������'\���d�,���p�:L��}<����)��H%X