BZh91AY&SYҦļ �_�Py����߰����P�=���ۜ�,vВ)�S���M&��mCjz��=@4���h�4Q�Q� =@  � $D�&CT�O4��O)�=M�6���b��M2dɈ��	�����$�&56���OS�hi�   5螺��(@@ �����)�M?R��%|`X4�i�� d��vp�BYf@m����~^c�ў~�we�ַ�",�zn~�,��}q�9S�T����gf�7	�)��ܙ��7���IF������e�^ѭ��N �dNI ���	L���r+9�o���5�z}�/��FH�&�vcWZ�m��^���V�s��5��fT�P��/�U�X�W���|s5I��ei���U��F89�Y���n
�5�H�Fs���P�S����3T�5Ta�I^��p�pJ�&Y�P'�.��_��֝֟�µ�u���bw�sy;�&�����l"-هJ��Qô�#�"̗�e8�^�-c�0&�=CaHfpL��d��MB�YQ90�R�t�_�4#k;Y��}���Fs�1��g)"��vo]��=O��V�u/�ҕ��J��e���VF�~����JA62.]?�ݶc$j+3�>+?){d[�}��t3$���x��[���T����NwZ&Gq-��c	H����23>D����bR�������d١���U�e�CD�'�RIUq��0��+X܆t����f0�-�H=i�j�&z��F�2���%�4f�DgΖ�q�c�ĽtR��N6;<J�G�ɳ],S�$�뤑P���9�P�&�ӣ�NDFܷ���8���=�ťl8��lm�q����P�ʮ��*�Bnh���g����d�Yc��c(��&�_!,W,��^ �@�&䤓L��и�Ф���G�	�g�- �-j�8�	Nl��ĵs�R
���k�WQ�˴�Ȑf-��s��g?�I��`�>X\M�i)U�}�0kY�8F�Vd�w�N^��3�����Q�i��7�m
t_Eh��
D��fR�ID�a���2өbb�c_"
}P�A1`��+�%�TpJ���w�T,!c�0��Q	����T:��=D���RD]j�@�b�aaf��ا.0��"2�u�E���	�p�[,�j��rr
���Iz��w$S�	*lK�