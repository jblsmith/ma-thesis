BZh91AY&SY� _�Py����߰����`�x�5�5j(   q�&LF& L�&@F �*`L�S@  �    dɓ��&	�F�!�I�H�OSj�4��h4= 4���q�&LF& L�&@F � �$	�&�Ai��S����M<���z���A��.X��O��,j|I��3h��Fk!#,�g�����2Ą�b2p���&u]:&ߨϲg��meZ���^�o���b����23+��h�4v�7���#�0���LB�8��<;p��w�Nj�G8�Vd���&޳��h��"�Y����"�����;� 23t���KF����Zv�^޻sS&�?"l0��_1��BMF��=�c>;�U'v�ƣ���H��`ž3��K�F��v�5�I����W�/e.SL����ݥ��V:0�;��p��mac<�c�&`T�Nt�nʢ6˶M�ѳę�ΰ���T�!9��dB�k���У��e�`JB��r��ɭ�l��+-�]�p����1�q��Ö͆�`֊I��R�ڣd�%�ZD!���.� z�J� h�k2͐$�>�iֲ8��J�qMB6���jZq%16����9�tC��1��MV6�&�7K�$
!
�]"#���0�\���L��Mr�Ή�)�Eu*�D$�	s�`�v'�|1$
�Uv$L8����v�R��B�P���C"}
��j�0��U�*jRZ�#��A��,ZB�`Ҽ��I�����3'�I3'NɅr|�S����N�E87�{O2��ܰ��n��ɵ�\�>s�n�,�]��\O���y�__ݪ��5���.v���,��2��Ok������gI��?I���z�S��[�xL�!'AQ*�)L�M.f���a"�1s,��i{������b�U���OL�5^)�Ӄ�:Lݓs�sT�X��8N�NUL�ͱ,YGɉ�y�e�Ɛ�z[[l�S.��:���7�]RѺ�
���\�J�8�DƐ���T���5Q쨳Lw35K�G�*�&G�21o�v#����ʔ�2bͷ�d�F���НM��-�NWV:%�D��Nق�֫Ψ���s�ɚt8ъ͙ܿ�\�T}�n�9'�����b�29�����8���n70l8�M�3b�R��B�x����a����h�;(C�z�0ر;����80�L�猳(o]'����`�)�]�t�P�KG�l�G����LY�,�b�*~�&7H�_�Y�%��k�.b�����ZK�x�>������s9�&��b;����;W��׋�ۻ�}�pr�tʡ��J~'l�2k�/T�INu�$;
/U����-N�+3�ɩ�i������<m��(�,�Ν�I����}�E��=΃���]&�Mn��%�R�ݬ�6��X2u���bjǽm��d�nl.�U)��r#�E�b��rl�͚kq�ͥrܺ#f�-=�	� �Oz�[�����o�mT��ڜm�����N��_�˝������QD�j��ݫ/�.�p� �8.