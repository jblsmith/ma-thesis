BZh91AY&SYN��� �_�py����߰����`���yǦ������`ڒ��#�ڀ�y  ��#@�  D��M      q�&�a22bh�A�L D�*�        �B�SOJ���A���  �SOS@�"iOE<���6 ��=OM'�4� �i�APT�����,�$����!U,�(>�?�h�"�(A,1D��!�KQx��2�P�QU�rA��vD���M'O!��Ws�[�֨�~�	��H�Sb�U0��S2�>�:�kH�J��I�R%(���{�OT�F��P����3��4�R�ln����a��[
��	J)TLɆev�P��*R�wQ	#�d�v����$&���2ˇ�#��c�z鬩E�6��}Ʒ3M����-3���_�"��8��',�j���s��ʤk�$Ϊ��K�y*�#�����lN��z&�MƳ�N���,e���ڝ!�)�eO�^e۰I�:3|��9��ӓ�fE��3������$R���	fd�t�^��"<9"=��d�:�5�!KQ�����/E@��eR��
����% ��Ř��/';��Q�b5g4u�m�F��Ѝ͡cCW���&�U䜁)$���,�A��0�k,�rђ�[%j ���dN�́F��g
� SB�r�.�+$#a�w@��I�$&mEAQ���E���@�sE�L�-8�e�Is�*�r�F$#���Ѳ�-+�2qF��X���FFbی٭Ըp�D8��tk9:�Ë�ٚi��|h��  {vF��$�I ��E=��jY����5U7aft�F��H�Ts��T/A�V�Bڭ!��|X!���F@�dMll�^�YWy�����;��ΌKG'�6ǌ`
m����UhuRǉK%�����Y�96G�ޘ��3�M$z%$)���%�~?_�Ȯ�cQ�2$���_�Fc�i����-è������M��v>t����~�C����"r�
I}���p��x>SMj�E.P�!�Y��*��*���Ap/X�_�>�;�^����4:F��׍&Wi��sAsRon������ӻ�i�u�h�
���s6�׎<G4��ͣ8	��Ǜ9?U� AX�pi#}�>�s���<��)�������0�����0��N��;C3��f�p��m:���?/-�7����P@D�,\��Ժd�l�j|agL^��=�g���')߼R�"꜉"�ʈ�J@b���>XG~�����0�s����iR=-k�tƉ��́�ʑ����:������g�p��hI���fM���*��u��3����/�����P����CId#�i9��7�K��r3l^5v�CgZ.�9�%��������!���J���9ћ;=� �v������E:Nġ5���wΎ0�:�X>���Ψ �FRN�炧j@͉'e��w$���s�E�[���)zu7&)V$I�ukvZ ��E.Z����w3ϙ�K�����
!�����!�:����¸7�`�YCPD�x�B�G��nWs������,� �����%��+В5��V�U�(:�JY�ΆB�aǳ�yr	,���ª�3�G�x��α��с��?����w$S�	�olp