BZh91AY&SY�c�� �߀Py����߰����P�lڣ��:����0I
zzBy)�	�m��M!�1#LA(A��MMGꙨh2 �� �I��
i�F����C�  �*�z4 �f�h2bi�� DMS�Oi6��L����P�  0H�5�"VB �I�����"�3�C����v��-�җ��qR����ё!D@BPr�j�f\\F������:�1��[�㍍d�*bx_��E �/"<�Zffd��r���?*���I#���V�b�DU��f[2s���� %(p�ik�S��q�9�ш8����{�����# �&���ش&�gj��"�k�Cغ��#%��ͦn��to���˙C@��#��f�wi�}
+����w�&�cg_>����ӽ3��5)�J-k;ѻN�4���5�UQ�剱4��X�S JE���h�6r�k�<�Yi�4袨���{8!m:�!!%��H �W&n8����ı),�����͂F�C���RM�`5���G��)(q*��qA6Pe-�1�d��\-s���S�Yg0��z<� 
�v-ү.�ź�h ����(���S�|�|�y($�q�:�����@kL�@�}���� ��-��s��K���4!� ��3	���-�%͢��*>�iT�<L��aqD~I�������J�w���h.$vX�р�َB~l�q����X�~<�1�=��>Η	�0�JZnNf�T����d��r��(��;�i�7�`>H�G��)A���b����E㓮/(��+�ʎ.K5%�821m �j4�r|�|��RR%~Q���'vL��5E�(p7��E�N6�]R�2�/R��U
�1�F�)p5T�� ���r[��t�J��2�X5�M�%cI��IJ�l�&A	0Xï�R`q�I,"q�%�i��c�PR�H�F���ܩ�(����0* X�t�Z!��Jpր�J-10���Is�58h��0�+)�lI��E��[Ja�8����F�UU0�b}Z��OȜ�:���H\��,�_��Z��Wj�,����dA�RH�g�|�[rQL�|�R��6E�E^Nu+*����5� ��0B�k��S1�b��i�+�5!��*�!q���=�N1�'!�8��ͫ2a��
��]up�̬RM��A�s��ɐg����w$S�	V;�0