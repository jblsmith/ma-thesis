BZh91AY&SY���b �_�Py����߰����`_3X Td  %	M��CD�����44M!��$�&�6�L0�0�4�2d�b`ɂd ф``8ɓ&# &L �# C�L�1�2`� 4a��!=E?D�&��y5=& �����\���$b�K�I-$&r~�H��U��O�ژ>�2�.�<�B��y?�d���	#d�dL�)KTz�Dʍk�l�s	f����ٜ*Ğ�N��uZ�uG��$��ZS��ػ�p�C�w�^�?y��J�����������Q�\���E$�A�SG����(��E���e���
&hQnZ(�F�����ކ�Un��Վ��bf�|��b���v^W#r��ld�nhcW�$1�^@x���S�LF3$��P.�ʓ��C#X%E$�TT�1��e��`S�V�۵�A�˻�� q�G4�sE���b� �AF�6?	�6+!
�k[ q�J�n(s�D��Yjq�!	����:*����;��9{"!K62�m�@��
��٨�Y�ҨQ�4*�(^6TE���D�8�A'6�6X�
c���V���3
���-�ƜkkE0]��䊊X��C�82�+n��%���b�$��\�$�H90L
lٖ*�l�AKd�t�$�D��0Kшⴎ4Q�b�AlRt\r�F���p����r8��r8�@�aأ\����ĝn���O��<JU)U󪪪���,�������阐�Q#>��R��8�xTB�;��zYT�e"��J�VW/-V�0�-(R���y^%,I{Y�b˫Zɒ����f�t�n���h.\�7�#�,�M��� �0h�2Pg����y��j,$q,A�7Kw#�J7Qb���W&"dQ����r�f{�ݛ=͑�J�R���$2���O㟬��S�y�ꓽ����-)B���H�ͳƱ�x�oG�2����n���0t�����G�ܒ?F�����r7�i/bx��w��L��H���:]��:R�=̀a7"����l>C��^��U�@ꌄ�J1^�o��)Q8J��T%��Т��Q�͑�k9&�ޔ�R!V����S3&��ђ�|]-|ҥ7L�5�r��Ծ��'���\���D�I!��<-Xb�ݹt��mg�%���&s	?V��$��8�wSS��3;Jr��ZV����Ÿ�Im��V��/���1W�y�=OL��mZ6�5GbH{��7,N��zoFkR���]K(s/'��	�S��2YB�o�d^I"��Z>��R>L"t�d��텊X��X�e�M3�1f�
[�d��2<LP�
֝����%v��.	!�b2�g+|0_S��>�~O)��_D�ln,9?}�'S�n�T?ds����y�ͥH͂�$�����pґ^b�*�ߨw:�B���ɲVm����Tv25�h�R��e�vosL[qMXLo�3�������;J�\3��&�,#�Fɸ�*g�7kL�S�/���ͯ���aªS���F�K&�M�(�۵��4pjku-���۪KC/��<̹����j�{�޾>�M�����1S2�n�G��$8�c����m�&����)�|��