BZh91AY&SY�M�? �߀Py����߰����`�O��/[�yY� JjJx�z#�i��2d�=54�h����=�?T        �S�j� �h     $��(ڙ��F�dz��CA�2=CM2d�L&F@��M#4i���z��5��Lj1 �,��j�ȃd(T1_���W~��o�j���똑��,��TF8LMW�5Y˅�As�G0���	5��q^�ϟ�kFq�P�rmP��B�Z�RV6$��D�PR�q�� ����a��Ϡd�I٦O�!qKzY6"G�*��+�c�q�F��XiL���a��$�S ��qC���(�!$�+B$���n�I��.�&��5�̆�=!�n����26L0�CN~�<����r1�ׁ���u��tP1鱲փZ^V�t�p��jÃ-N�s�JZ��N�1�w�	�?�qy��,b&\�m_|{󊻡}��{�SmBd��1�B��*9Q�wE�*��8P�n�+��N�Jgt��	���b��zaH"���d\P*�Z�X��sl�+fЁ� 9�;`ta�Khx��N|j#BX@����V*IB�X%!�Lh�f�Ce�Q[	�."���ZV�lc�
bO?Q�8��l���HBNI$�Th��)�6s3�b��9��UR%_CTi]t Z ��"Q#!�/bZ^�b$#�"S��%A���	�UI��$N	��TcNUEO����P�&j��`�j��4i�aY3O�F�Q�f1 ��Y�Q��e�Z�O �u|��D|L4�)�v����]2z��HBRRvf0od~� ���뮳rB":J!��u8��z�n#F���"9�q48�p4m��D��݇��D{��P���rE�c.JP�Cq��ı�Д&( 7V!��=& �h+X/1-�7�<(�x�0��̙&��;����"c��+0J�P0jS������̰b��?D!8��g�Ղ��:�T`��a~i�d�T�ˡXTEĴ�aq=���v�,k9W`@4!L�� �0�:��<����7p	��`�_ɦ,���r0�q4X5���9:�a$�_��z
��!`d1���.-?�aA�JS^�� �`v�HԻ.��@^��w� ��9��&J��������I.ҥCNO�,H`Ld������:�E9�GE��f���Pw���b�(I�Bĉ�&H $T�4T<�D	@L����q|�FA�ڄ.e �:H$J�i1|���cذ�	xLJ����y�w��� 0���15��&R�b#�Z6I�`0��:�Q�P�2�������m0���_�
5�AGJ�1p���J���_a�7��\5��m?1_Ț3�,�EYj3'q`*��24���B��t)mm2���f5�k�Y�y���^`n#]�W%0+�Tz@���k��F�7f��L�t#R���&��:�u���́.����c�CV6��ܑN$+�l�